
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library ieee_proposed;
use ieee_proposed.fixed_pkg.all;


-- Positive half of the sigmoid function
entity sigmoid is
port (
    clk: in std_logic;
    rst: in std_logic;
    datain: in std_logic_vector (16 - 2 downto 0);
    validin: in std_logic;
    dataout: out std_logic_vector (16 - 2 downto 0);
    validout: out std_logic);
end sigmoid;

architecture Behavioural of sigmoid is

constant PIPE_LEN: natural := 630;

signal pipe_in: std_logic_vector (PIPE_LEN - 1 downto 0);
signal pipe_out: std_logic_vector (PIPE_LEN - 1 downto 0);

begin

process (clk, rst) is
begin
    if (rising_edge(clk)) then
        if (rst = '0') then
            pipe_out <= (others => '0');
        else
            pipe_out <= pipe_in;
        end if;
    end if;
end process;

-- data is present a cycle later
process (clk, rst) is
begin
    if (rising_edge(clk)) then
        if (rst = '0') then
            validout <= '0';
        else
            validout <= validin;
        end if;
    end if;
end process;

-- auto-generated combinational code starts here
pipe_in (0) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (1) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (2) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (3) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (4) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (5) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (6) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (7) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (8) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (9) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (10) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (11) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (12) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (13) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (14) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (15) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (16) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (17) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (18) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (19) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (20) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (21) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (22) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (23) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (24) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (25) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (26) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (27) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (28) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (29) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (30) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (31) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (32) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (33) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (34) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (35) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (36) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (37) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (38) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (39) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (40) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (41) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (42) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (43) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (44) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (45) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (46) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (47) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (48) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (49) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (50) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (51) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (52) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (53) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (54) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (55) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (56) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (57) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (58) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (59) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (60) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (61) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (62) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (63) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (64) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (65) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (66) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (67) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (68) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (69) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (70) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (71) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (72) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (73) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (74) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (75) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (76) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (77) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (78) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (79) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (80) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (81) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (82) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (83) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (84) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (85) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (86) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (87) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (88) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (89) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (90) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (91) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (92) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (93) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (94) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (95) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (96) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (97) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (98) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (99) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (100) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (101) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (102) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (103) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and datain (7) = '1' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (104) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (105) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (106) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (107) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (108) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (109) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (110) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (111) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (112) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (113) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (114) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (115) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (116) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (117) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (118) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (119) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (120) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (121) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (122) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (123) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (124) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (125) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (126) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (127) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (128) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (129) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (130) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and (true) else '0';
pipe_in (131) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and (true) else '0';
pipe_in (132) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and datain (7) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (133) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (134) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and (true) else '0';
pipe_in (135) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and (true) else '0';
pipe_in (136) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (9) = '1' and (true) else '0';
pipe_in (137) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (11) = '1' and (true) else '0';
pipe_in (138) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '1' and (true) else '0';
dataout (0) <= '1' when pipe_out (0) = '1' or pipe_out (1) = '1' or pipe_out (2) = '1' or pipe_out (3) = '1' or pipe_out (4) = '1' or pipe_out (5) = '1' or pipe_out (6) = '1' or pipe_out (7) = '1' or pipe_out (8) = '1' or pipe_out (9) = '1' or pipe_out (10) = '1' or pipe_out (11) = '1' or pipe_out (12) = '1' or pipe_out (13) = '1' or pipe_out (14) = '1' or pipe_out (15) = '1' or pipe_out (16) = '1' or pipe_out (17) = '1' or pipe_out (18) = '1' or pipe_out (19) = '1' or pipe_out (20) = '1' or pipe_out (21) = '1' or pipe_out (22) = '1' or pipe_out (23) = '1' or pipe_out (24) = '1' or pipe_out (25) = '1' or pipe_out (26) = '1' or pipe_out (27) = '1' or pipe_out (28) = '1' or pipe_out (29) = '1' or pipe_out (30) = '1' or pipe_out (31) = '1' or pipe_out (32) = '1' or pipe_out (33) = '1' or pipe_out (34) = '1' or pipe_out (35) = '1' or pipe_out (36) = '1' or pipe_out (37) = '1' or pipe_out (38) = '1' or pipe_out (39) = '1' or pipe_out (40) = '1' or pipe_out (41) = '1' or pipe_out (42) = '1' or pipe_out (43) = '1' or pipe_out (44) = '1' or pipe_out (45) = '1' or pipe_out (46) = '1' or pipe_out (47) = '1' or pipe_out (48) = '1' or pipe_out (49) = '1' or pipe_out (50) = '1' or pipe_out (51) = '1' or pipe_out (52) = '1' or pipe_out (53) = '1' or pipe_out (54) = '1' or pipe_out (55) = '1' or pipe_out (56) = '1' or pipe_out (57) = '1' or pipe_out (58) = '1' or pipe_out (59) = '1' or pipe_out (60) = '1' or pipe_out (61) = '1' or pipe_out (62) = '1' or pipe_out (63) = '1' or pipe_out (64) = '1' or pipe_out (65) = '1' or pipe_out (66) = '1' or pipe_out (67) = '1' or pipe_out (68) = '1' or pipe_out (69) = '1' or pipe_out (70) = '1' or pipe_out (71) = '1' or pipe_out (72) = '1' or pipe_out (73) = '1' or pipe_out (74) = '1' or pipe_out (75) = '1' or pipe_out (76) = '1' or pipe_out (77) = '1' or pipe_out (78) = '1' or pipe_out (79) = '1' or pipe_out (80) = '1' or pipe_out (81) = '1' or pipe_out (82) = '1' or pipe_out (83) = '1' or pipe_out (84) = '1' or pipe_out (85) = '1' or pipe_out (86) = '1' or pipe_out (87) = '1' or pipe_out (88) = '1' or pipe_out (89) = '1' or pipe_out (90) = '1' or pipe_out (91) = '1' or pipe_out (92) = '1' or pipe_out (93) = '1' or pipe_out (94) = '1' or pipe_out (95) = '1' or pipe_out (96) = '1' or pipe_out (97) = '1' or pipe_out (98) = '1' or pipe_out (99) = '1' or pipe_out (100) = '1' or pipe_out (101) = '1' or pipe_out (102) = '1' or pipe_out (103) = '1' or pipe_out (104) = '1' or pipe_out (105) = '1' or pipe_out (106) = '1' or pipe_out (107) = '1' or pipe_out (108) = '1' or pipe_out (109) = '1' or pipe_out (110) = '1' or pipe_out (111) = '1' or pipe_out (112) = '1' or pipe_out (113) = '1' or pipe_out (114) = '1' or pipe_out (115) = '1' or pipe_out (116) = '1' or pipe_out (117) = '1' or pipe_out (118) = '1' or pipe_out (119) = '1' or pipe_out (120) = '1' or pipe_out (121) = '1' or pipe_out (122) = '1' or pipe_out (123) = '1' or pipe_out (124) = '1' or pipe_out (125) = '1' or pipe_out (126) = '1' or pipe_out (127) = '1' or pipe_out (128) = '1' or pipe_out (129) = '1' or pipe_out (130) = '1' or pipe_out (131) = '1' or pipe_out (132) = '1' or pipe_out (133) = '1' or pipe_out (134) = '1' or pipe_out (135) = '1' or pipe_out (136) = '1' or pipe_out (137) = '1' or pipe_out (138) = '1' or (false) else '0';
pipe_in (139) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (140) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (141) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (142) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (143) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (144) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (145) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (146) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (147) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (148) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (149) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (150) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (151) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (152) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (153) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (154) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (155) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (156) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (157) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (158) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (159) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (160) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (161) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (162) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (163) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '1' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (164) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (165) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (166) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (167) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (168) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (169) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (170) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (171) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (172) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (173) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (174) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (175) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (176) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (177) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (178) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (179) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (180) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (181) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (182) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (183) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (184) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (185) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (186) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (187) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (188) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (189) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (190) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (191) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (192) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (193) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (3) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (194) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (195) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (196) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (3) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (197) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (4) = '0' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (198) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (199) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (200) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (201) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (202) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (203) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (204) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (205) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (206) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (207) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (208) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (209) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (210) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (211) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (212) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (213) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (214) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (215) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (216) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (217) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (218) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (219) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (220) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (221) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (222) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (223) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (224) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (225) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (226) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (227) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (228) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (229) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (230) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (231) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (232) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (233) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (234) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (235) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and (true) else '0';
pipe_in (236) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and (true) else '0';
pipe_in (237) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (238) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and (true) else '0';
pipe_in (239) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (240) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and (true) else '0';
pipe_in (241) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (242) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (243) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and (true) else '0';
pipe_in (244) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (9) = '1' and (true) else '0';
pipe_in (245) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and (true) else '0';
pipe_in (246) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (11) = '1' and (true) else '0';
pipe_in (247) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '1' and (true) else '0';
dataout (1) <= '1' when pipe_out (139) = '1' or pipe_out (140) = '1' or pipe_out (141) = '1' or pipe_out (142) = '1' or pipe_out (143) = '1' or pipe_out (144) = '1' or pipe_out (145) = '1' or pipe_out (146) = '1' or pipe_out (147) = '1' or pipe_out (148) = '1' or pipe_out (149) = '1' or pipe_out (150) = '1' or pipe_out (151) = '1' or pipe_out (152) = '1' or pipe_out (153) = '1' or pipe_out (154) = '1' or pipe_out (155) = '1' or pipe_out (156) = '1' or pipe_out (157) = '1' or pipe_out (158) = '1' or pipe_out (159) = '1' or pipe_out (160) = '1' or pipe_out (161) = '1' or pipe_out (162) = '1' or pipe_out (163) = '1' or pipe_out (164) = '1' or pipe_out (165) = '1' or pipe_out (166) = '1' or pipe_out (167) = '1' or pipe_out (168) = '1' or pipe_out (169) = '1' or pipe_out (170) = '1' or pipe_out (171) = '1' or pipe_out (172) = '1' or pipe_out (173) = '1' or pipe_out (174) = '1' or pipe_out (175) = '1' or pipe_out (176) = '1' or pipe_out (177) = '1' or pipe_out (178) = '1' or pipe_out (179) = '1' or pipe_out (180) = '1' or pipe_out (181) = '1' or pipe_out (182) = '1' or pipe_out (183) = '1' or pipe_out (184) = '1' or pipe_out (185) = '1' or pipe_out (186) = '1' or pipe_out (187) = '1' or pipe_out (188) = '1' or pipe_out (189) = '1' or pipe_out (190) = '1' or pipe_out (191) = '1' or pipe_out (192) = '1' or pipe_out (193) = '1' or pipe_out (194) = '1' or pipe_out (195) = '1' or pipe_out (196) = '1' or pipe_out (197) = '1' or pipe_out (198) = '1' or pipe_out (199) = '1' or pipe_out (200) = '1' or pipe_out (201) = '1' or pipe_out (202) = '1' or pipe_out (203) = '1' or pipe_out (204) = '1' or pipe_out (205) = '1' or pipe_out (206) = '1' or pipe_out (207) = '1' or pipe_out (208) = '1' or pipe_out (209) = '1' or pipe_out (210) = '1' or pipe_out (211) = '1' or pipe_out (212) = '1' or pipe_out (213) = '1' or pipe_out (214) = '1' or pipe_out (215) = '1' or pipe_out (216) = '1' or pipe_out (217) = '1' or pipe_out (218) = '1' or pipe_out (219) = '1' or pipe_out (220) = '1' or pipe_out (221) = '1' or pipe_out (222) = '1' or pipe_out (223) = '1' or pipe_out (224) = '1' or pipe_out (225) = '1' or pipe_out (226) = '1' or pipe_out (227) = '1' or pipe_out (228) = '1' or pipe_out (229) = '1' or pipe_out (230) = '1' or pipe_out (231) = '1' or pipe_out (232) = '1' or pipe_out (233) = '1' or pipe_out (234) = '1' or pipe_out (235) = '1' or pipe_out (236) = '1' or pipe_out (237) = '1' or pipe_out (238) = '1' or pipe_out (239) = '1' or pipe_out (240) = '1' or pipe_out (241) = '1' or pipe_out (242) = '1' or pipe_out (243) = '1' or pipe_out (244) = '1' or pipe_out (245) = '1' or pipe_out (246) = '1' or pipe_out (247) = '1' or (false) else '0';
pipe_in (248) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (249) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (250) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (251) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (252) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (253) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (254) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (255) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (256) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (257) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (258) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (259) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (260) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (261) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (262) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (263) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (264) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (265) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (266) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (267) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (268) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (269) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (270) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (271) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (272) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (273) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (274) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (275) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (276) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (277) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (278) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (4) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (279) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (280) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (281) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (282) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (283) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (284) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (285) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (286) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (287) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (288) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (289) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (290) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (291) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (292) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (293) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (294) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (295) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (296) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (297) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (298) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (299) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (300) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (301) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (302) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and (true) else '0';
pipe_in (303) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (304) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (305) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (306) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (307) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (308) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (309) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (310) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (311) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and (true) else '0';
pipe_in (312) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and (true) else '0';
pipe_in (313) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (314) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and (true) else '0';
pipe_in (315) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (316) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (9) = '1' and (true) else '0';
pipe_in (317) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (318) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and (true) else '0';
pipe_in (319) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (11) = '1' and (true) else '0';
pipe_in (320) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '1' and (true) else '0';
dataout (2) <= '1' when pipe_out (248) = '1' or pipe_out (249) = '1' or pipe_out (250) = '1' or pipe_out (251) = '1' or pipe_out (252) = '1' or pipe_out (253) = '1' or pipe_out (254) = '1' or pipe_out (255) = '1' or pipe_out (256) = '1' or pipe_out (257) = '1' or pipe_out (258) = '1' or pipe_out (259) = '1' or pipe_out (260) = '1' or pipe_out (261) = '1' or pipe_out (262) = '1' or pipe_out (263) = '1' or pipe_out (264) = '1' or pipe_out (265) = '1' or pipe_out (266) = '1' or pipe_out (267) = '1' or pipe_out (268) = '1' or pipe_out (269) = '1' or pipe_out (270) = '1' or pipe_out (271) = '1' or pipe_out (272) = '1' or pipe_out (273) = '1' or pipe_out (274) = '1' or pipe_out (275) = '1' or pipe_out (276) = '1' or pipe_out (277) = '1' or pipe_out (278) = '1' or pipe_out (279) = '1' or pipe_out (280) = '1' or pipe_out (281) = '1' or pipe_out (282) = '1' or pipe_out (283) = '1' or pipe_out (284) = '1' or pipe_out (285) = '1' or pipe_out (286) = '1' or pipe_out (287) = '1' or pipe_out (288) = '1' or pipe_out (289) = '1' or pipe_out (290) = '1' or pipe_out (291) = '1' or pipe_out (292) = '1' or pipe_out (293) = '1' or pipe_out (294) = '1' or pipe_out (295) = '1' or pipe_out (296) = '1' or pipe_out (297) = '1' or pipe_out (298) = '1' or pipe_out (299) = '1' or pipe_out (300) = '1' or pipe_out (301) = '1' or pipe_out (302) = '1' or pipe_out (303) = '1' or pipe_out (304) = '1' or pipe_out (305) = '1' or pipe_out (306) = '1' or pipe_out (307) = '1' or pipe_out (308) = '1' or pipe_out (309) = '1' or pipe_out (310) = '1' or pipe_out (311) = '1' or pipe_out (312) = '1' or pipe_out (313) = '1' or pipe_out (314) = '1' or pipe_out (315) = '1' or pipe_out (316) = '1' or pipe_out (317) = '1' or pipe_out (318) = '1' or pipe_out (319) = '1' or pipe_out (320) = '1' or (false) else '0';
pipe_in (321) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (322) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (323) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (324) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (325) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (326) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (327) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (328) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (329) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (330) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (331) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (332) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (333) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (334) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (335) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (336) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (337) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (338) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (339) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (340) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (341) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (342) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (343) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (344) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (345) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (346) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (347) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (348) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (349) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (350) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (351) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (352) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (353) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (354) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (355) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (356) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (357) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (358) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (359) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (360) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (361) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (362) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (363) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (364) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (365) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (366) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (367) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (368) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (369) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (370) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (371) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (372) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (373) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (374) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (375) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (376) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (377) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and (true) else '0';
pipe_in (378) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (379) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (380) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (381) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (382) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (383) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (384) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and (true) else '0';
pipe_in (385) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and (true) else '0';
pipe_in (386) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and (true) else '0';
pipe_in (387) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (388) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (9) = '1' and (true) else '0';
pipe_in (389) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (390) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and (true) else '0';
pipe_in (391) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (11) = '1' and (true) else '0';
pipe_in (392) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '1' and (true) else '0';
dataout (3) <= '1' when pipe_out (321) = '1' or pipe_out (322) = '1' or pipe_out (323) = '1' or pipe_out (324) = '1' or pipe_out (325) = '1' or pipe_out (326) = '1' or pipe_out (327) = '1' or pipe_out (328) = '1' or pipe_out (329) = '1' or pipe_out (330) = '1' or pipe_out (331) = '1' or pipe_out (332) = '1' or pipe_out (333) = '1' or pipe_out (334) = '1' or pipe_out (335) = '1' or pipe_out (336) = '1' or pipe_out (337) = '1' or pipe_out (338) = '1' or pipe_out (339) = '1' or pipe_out (340) = '1' or pipe_out (341) = '1' or pipe_out (342) = '1' or pipe_out (343) = '1' or pipe_out (344) = '1' or pipe_out (345) = '1' or pipe_out (346) = '1' or pipe_out (347) = '1' or pipe_out (348) = '1' or pipe_out (349) = '1' or pipe_out (350) = '1' or pipe_out (351) = '1' or pipe_out (352) = '1' or pipe_out (353) = '1' or pipe_out (354) = '1' or pipe_out (355) = '1' or pipe_out (356) = '1' or pipe_out (357) = '1' or pipe_out (358) = '1' or pipe_out (359) = '1' or pipe_out (360) = '1' or pipe_out (361) = '1' or pipe_out (362) = '1' or pipe_out (363) = '1' or pipe_out (364) = '1' or pipe_out (365) = '1' or pipe_out (366) = '1' or pipe_out (367) = '1' or pipe_out (368) = '1' or pipe_out (369) = '1' or pipe_out (370) = '1' or pipe_out (371) = '1' or pipe_out (372) = '1' or pipe_out (373) = '1' or pipe_out (374) = '1' or pipe_out (375) = '1' or pipe_out (376) = '1' or pipe_out (377) = '1' or pipe_out (378) = '1' or pipe_out (379) = '1' or pipe_out (380) = '1' or pipe_out (381) = '1' or pipe_out (382) = '1' or pipe_out (383) = '1' or pipe_out (384) = '1' or pipe_out (385) = '1' or pipe_out (386) = '1' or pipe_out (387) = '1' or pipe_out (388) = '1' or pipe_out (389) = '1' or pipe_out (390) = '1' or pipe_out (391) = '1' or pipe_out (392) = '1' or (false) else '0';
pipe_in (393) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (394) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (395) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (396) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (397) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (398) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (399) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (400) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (401) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (402) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (403) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (404) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (405) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (406) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (407) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (408) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (409) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (410) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (411) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (412) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (413) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (414) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (415) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (416) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (417) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (418) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (419) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (420) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (421) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (422) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (423) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (424) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (425) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (426) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (427) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (428) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (429) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (430) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (431) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (432) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (433) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (434) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (435) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (436) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (437) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (438) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (439) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (440) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (441) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (442) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (443) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and (true) else '0';
pipe_in (444) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (445) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (446) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (447) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (448) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (449) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (450) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (451) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (452) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (453) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (454) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (455) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (456) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (457) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and (true) else '0';
pipe_in (458) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (459) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (460) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and (true) else '0';
pipe_in (461) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and (true) else '0';
pipe_in (462) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (463) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (464) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and (true) else '0';
pipe_in (465) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (11) = '1' and (true) else '0';
pipe_in (466) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '1' and (true) else '0';
dataout (4) <= '1' when pipe_out (393) = '1' or pipe_out (394) = '1' or pipe_out (395) = '1' or pipe_out (396) = '1' or pipe_out (397) = '1' or pipe_out (398) = '1' or pipe_out (399) = '1' or pipe_out (400) = '1' or pipe_out (401) = '1' or pipe_out (402) = '1' or pipe_out (403) = '1' or pipe_out (404) = '1' or pipe_out (405) = '1' or pipe_out (406) = '1' or pipe_out (407) = '1' or pipe_out (408) = '1' or pipe_out (409) = '1' or pipe_out (410) = '1' or pipe_out (411) = '1' or pipe_out (412) = '1' or pipe_out (413) = '1' or pipe_out (414) = '1' or pipe_out (415) = '1' or pipe_out (416) = '1' or pipe_out (417) = '1' or pipe_out (418) = '1' or pipe_out (419) = '1' or pipe_out (420) = '1' or pipe_out (421) = '1' or pipe_out (422) = '1' or pipe_out (423) = '1' or pipe_out (424) = '1' or pipe_out (425) = '1' or pipe_out (426) = '1' or pipe_out (427) = '1' or pipe_out (428) = '1' or pipe_out (429) = '1' or pipe_out (430) = '1' or pipe_out (431) = '1' or pipe_out (432) = '1' or pipe_out (433) = '1' or pipe_out (434) = '1' or pipe_out (435) = '1' or pipe_out (436) = '1' or pipe_out (437) = '1' or pipe_out (438) = '1' or pipe_out (439) = '1' or pipe_out (440) = '1' or pipe_out (441) = '1' or pipe_out (442) = '1' or pipe_out (443) = '1' or pipe_out (444) = '1' or pipe_out (445) = '1' or pipe_out (446) = '1' or pipe_out (447) = '1' or pipe_out (448) = '1' or pipe_out (449) = '1' or pipe_out (450) = '1' or pipe_out (451) = '1' or pipe_out (452) = '1' or pipe_out (453) = '1' or pipe_out (454) = '1' or pipe_out (455) = '1' or pipe_out (456) = '1' or pipe_out (457) = '1' or pipe_out (458) = '1' or pipe_out (459) = '1' or pipe_out (460) = '1' or pipe_out (461) = '1' or pipe_out (462) = '1' or pipe_out (463) = '1' or pipe_out (464) = '1' or pipe_out (465) = '1' or pipe_out (466) = '1' or (false) else '0';
pipe_in (467) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (468) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (469) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (470) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (471) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (472) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (473) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (474) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (475) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (476) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (477) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (478) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (479) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (480) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (481) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (482) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (483) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (484) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (485) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (486) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (487) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (488) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (489) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (490) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (491) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (492) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (493) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (494) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (495) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (496) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (497) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (498) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (499) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (500) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (501) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (502) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (503) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (504) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (505) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (506) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (507) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (508) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (509) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (510) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (511) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (512) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (513) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (514) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (515) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (516) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (517) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (518) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (519) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and (true) else '0';
pipe_in (520) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (521) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (522) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (523) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (524) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (525) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (526) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (527) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (528) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (529) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (530) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and (true) else '0';
pipe_in (531) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '0' and datain (7) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (532) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (533) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and (true) else '0';
pipe_in (534) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (535) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (536) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and (true) else '0';
pipe_in (537) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and (true) else '0';
pipe_in (538) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (539) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (540) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and (true) else '0';
pipe_in (541) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (11) = '1' and (true) else '0';
pipe_in (542) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '1' and (true) else '0';
dataout (5) <= '1' when pipe_out (467) = '1' or pipe_out (468) = '1' or pipe_out (469) = '1' or pipe_out (470) = '1' or pipe_out (471) = '1' or pipe_out (472) = '1' or pipe_out (473) = '1' or pipe_out (474) = '1' or pipe_out (475) = '1' or pipe_out (476) = '1' or pipe_out (477) = '1' or pipe_out (478) = '1' or pipe_out (479) = '1' or pipe_out (480) = '1' or pipe_out (481) = '1' or pipe_out (482) = '1' or pipe_out (483) = '1' or pipe_out (484) = '1' or pipe_out (485) = '1' or pipe_out (486) = '1' or pipe_out (487) = '1' or pipe_out (488) = '1' or pipe_out (489) = '1' or pipe_out (490) = '1' or pipe_out (491) = '1' or pipe_out (492) = '1' or pipe_out (493) = '1' or pipe_out (494) = '1' or pipe_out (495) = '1' or pipe_out (496) = '1' or pipe_out (497) = '1' or pipe_out (498) = '1' or pipe_out (499) = '1' or pipe_out (500) = '1' or pipe_out (501) = '1' or pipe_out (502) = '1' or pipe_out (503) = '1' or pipe_out (504) = '1' or pipe_out (505) = '1' or pipe_out (506) = '1' or pipe_out (507) = '1' or pipe_out (508) = '1' or pipe_out (509) = '1' or pipe_out (510) = '1' or pipe_out (511) = '1' or pipe_out (512) = '1' or pipe_out (513) = '1' or pipe_out (514) = '1' or pipe_out (515) = '1' or pipe_out (516) = '1' or pipe_out (517) = '1' or pipe_out (518) = '1' or pipe_out (519) = '1' or pipe_out (520) = '1' or pipe_out (521) = '1' or pipe_out (522) = '1' or pipe_out (523) = '1' or pipe_out (524) = '1' or pipe_out (525) = '1' or pipe_out (526) = '1' or pipe_out (527) = '1' or pipe_out (528) = '1' or pipe_out (529) = '1' or pipe_out (530) = '1' or pipe_out (531) = '1' or pipe_out (532) = '1' or pipe_out (533) = '1' or pipe_out (534) = '1' or pipe_out (535) = '1' or pipe_out (536) = '1' or pipe_out (537) = '1' or pipe_out (538) = '1' or pipe_out (539) = '1' or pipe_out (540) = '1' or pipe_out (541) = '1' or pipe_out (542) = '1' or (false) else '0';
pipe_in (543) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (544) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (545) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (546) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (547) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (548) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (549) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (550) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (551) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (552) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (553) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (554) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (555) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (556) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (557) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (558) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (559) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (560) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (561) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (562) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (563) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (564) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (565) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (566) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (567) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (568) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (569) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (570) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (571) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (572) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (573) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (574) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (575) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (576) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (577) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (578) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (579) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (580) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (581) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (582) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (583) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (584) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (585) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (586) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (587) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and (true) else '0';
pipe_in (588) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (589) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (590) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (591) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (592) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and (true) else '0';
pipe_in (593) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (594) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (595) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (596) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (597) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (598) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (599) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (600) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (601) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and (true) else '0';
pipe_in (602) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (603) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and (true) else '0';
pipe_in (604) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (605) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (606) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (8) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (607) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and (true) else '0';
pipe_in (608) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and (true) else '0';
pipe_in (609) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (610) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (611) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (10) = '1' and datain (8) = '1' and (true) else '0';
pipe_in (612) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (11) = '1' and (true) else '0';
pipe_in (613) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '1' and (true) else '0';
dataout (6) <= '1' when pipe_out (543) = '1' or pipe_out (544) = '1' or pipe_out (545) = '1' or pipe_out (546) = '1' or pipe_out (547) = '1' or pipe_out (548) = '1' or pipe_out (549) = '1' or pipe_out (550) = '1' or pipe_out (551) = '1' or pipe_out (552) = '1' or pipe_out (553) = '1' or pipe_out (554) = '1' or pipe_out (555) = '1' or pipe_out (556) = '1' or pipe_out (557) = '1' or pipe_out (558) = '1' or pipe_out (559) = '1' or pipe_out (560) = '1' or pipe_out (561) = '1' or pipe_out (562) = '1' or pipe_out (563) = '1' or pipe_out (564) = '1' or pipe_out (565) = '1' or pipe_out (566) = '1' or pipe_out (567) = '1' or pipe_out (568) = '1' or pipe_out (569) = '1' or pipe_out (570) = '1' or pipe_out (571) = '1' or pipe_out (572) = '1' or pipe_out (573) = '1' or pipe_out (574) = '1' or pipe_out (575) = '1' or pipe_out (576) = '1' or pipe_out (577) = '1' or pipe_out (578) = '1' or pipe_out (579) = '1' or pipe_out (580) = '1' or pipe_out (581) = '1' or pipe_out (582) = '1' or pipe_out (583) = '1' or pipe_out (584) = '1' or pipe_out (585) = '1' or pipe_out (586) = '1' or pipe_out (587) = '1' or pipe_out (588) = '1' or pipe_out (589) = '1' or pipe_out (590) = '1' or pipe_out (591) = '1' or pipe_out (592) = '1' or pipe_out (593) = '1' or pipe_out (594) = '1' or pipe_out (595) = '1' or pipe_out (596) = '1' or pipe_out (597) = '1' or pipe_out (598) = '1' or pipe_out (599) = '1' or pipe_out (600) = '1' or pipe_out (601) = '1' or pipe_out (602) = '1' or pipe_out (603) = '1' or pipe_out (604) = '1' or pipe_out (605) = '1' or pipe_out (606) = '1' or pipe_out (607) = '1' or pipe_out (608) = '1' or pipe_out (609) = '1' or pipe_out (610) = '1' or pipe_out (611) = '1' or pipe_out (612) = '1' or pipe_out (613) = '1' or (false) else '0';
pipe_in (614) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (615) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (616) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (617) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (618) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (619) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and (true) else '0';
pipe_in (620) <= '1' when datain (14) = '0' and datain (13) = '1' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and (true) else '0';
pipe_in (621) <= '1' when datain (14) = '0' and datain (13) = '0' and (true) else '0';
dataout (7) <= '1' when pipe_out (614) = '1' or pipe_out (615) = '1' or pipe_out (616) = '1' or pipe_out (617) = '1' or pipe_out (618) = '1' or pipe_out (619) = '1' or pipe_out (620) = '1' or pipe_out (621) = '1' or (false) else '0';
pipe_in (622) <= '1' when datain (13) = '1' and datain (10) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (623) <= '1' when datain (13) = '1' and datain (10) = '1' and datain (7) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (624) <= '1' when datain (13) = '1' and datain (10) = '1' and datain (7) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (625) <= '1' when datain (13) = '1' and datain (10) = '1' and datain (9) = '1' and (true) else '0';
pipe_in (626) <= '1' when datain (13) = '1' and datain (10) = '1' and datain (8) = '1' and (true) else '0';
pipe_in (627) <= '1' when datain (13) = '1' and datain (11) = '1' and (true) else '0';
pipe_in (628) <= '1' when datain (13) = '1' and datain (12) = '1' and (true) else '0';
pipe_in (629) <= '1' when datain (14) = '1' and (true) else '0';
dataout (8) <= '1' when pipe_out (622) = '1' or pipe_out (623) = '1' or pipe_out (624) = '1' or pipe_out (625) = '1' or pipe_out (626) = '1' or pipe_out (627) = '1' or pipe_out (628) = '1' or pipe_out (629) = '1' or (false) else '0';
dataout (9) <= '0';

dataout (10) <= '0';

dataout (11) <= '0';

dataout (12) <= '0';

dataout (13) <= '0';

dataout (14) <= '0';


end Behavioural;
