
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library ieee_proposed;
use ieee_proposed.fixed_pkg.all;


-- Positive half of the sigmoidgrad function
entity sigmoidgrad is
port (
    clk: in std_logic;
    rst: in std_logic;
    datain: in std_logic_vector (16 - 2 downto 0);
    validin: in std_logic;
    dataout: out std_logic_vector (16 - 2 downto 0);
    validout: out std_logic);
end sigmoidgrad;

architecture Behavioural of sigmoidgrad is

constant PIPE_LEN: natural := 296;

signal pipe_in: std_logic_vector (PIPE_LEN - 1 downto 0);
signal pipe_out: std_logic_vector (PIPE_LEN - 1 downto 0);

begin

process (clk, rst) is
begin
    if (rising_edge(clk)) then
        if (rst = '0') then
            pipe_out <= (others => '0');
        else
            pipe_out <= pipe_in;
        end if;
    end if;
end process;

-- data is present a cycle later
process (clk, rst) is
begin
    if (rising_edge(clk)) then
        if (rst = '0') then
            validout <= '0';
        else
            validout <= validin;
        end if;
    end if;
end process;

-- auto-generated combinational code starts here
pipe_in (0) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (1) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (2) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (3) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (4) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (5) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (6) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (7) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (8) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (9) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (10) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (11) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (12) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (13) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (14) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (15) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (16) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (17) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (18) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (19) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (20) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (21) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (22) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (23) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (24) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (25) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (26) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (27) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (28) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (29) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (30) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (31) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (32) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (33) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (34) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (4) = '0' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (35) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (36) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (37) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (38) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (39) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (40) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (41) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (42) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (43) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (44) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (45) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (46) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (47) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (48) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (49) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (50) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (51) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (52) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (53) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (54) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (55) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (56) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (3) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (57) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (58) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (59) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (60) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (61) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (62) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (63) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (64) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (65) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (66) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (67) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (68) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (69) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (70) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (71) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (72) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (73) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (74) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (75) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (76) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (77) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and (true) else '0';
pipe_in (78) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (79) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (80) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (81) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (82) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (83) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (84) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (85) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (86) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and (true) else '0';
pipe_in (87) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (88) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (89) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (90) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (91) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (92) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and (true) else '0';
pipe_in (93) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (94) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (95) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (96) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and (true) else '0';
pipe_in (97) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (98) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (0) = '1' and (true) else '0';
dataout (0) <= '1' when pipe_out (0) = '1' or pipe_out (1) = '1' or pipe_out (2) = '1' or pipe_out (3) = '1' or pipe_out (4) = '1' or pipe_out (5) = '1' or pipe_out (6) = '1' or pipe_out (7) = '1' or pipe_out (8) = '1' or pipe_out (9) = '1' or pipe_out (10) = '1' or pipe_out (11) = '1' or pipe_out (12) = '1' or pipe_out (13) = '1' or pipe_out (14) = '1' or pipe_out (15) = '1' or pipe_out (16) = '1' or pipe_out (17) = '1' or pipe_out (18) = '1' or pipe_out (19) = '1' or pipe_out (20) = '1' or pipe_out (21) = '1' or pipe_out (22) = '1' or pipe_out (23) = '1' or pipe_out (24) = '1' or pipe_out (25) = '1' or pipe_out (26) = '1' or pipe_out (27) = '1' or pipe_out (28) = '1' or pipe_out (29) = '1' or pipe_out (30) = '1' or pipe_out (31) = '1' or pipe_out (32) = '1' or pipe_out (33) = '1' or pipe_out (34) = '1' or pipe_out (35) = '1' or pipe_out (36) = '1' or pipe_out (37) = '1' or pipe_out (38) = '1' or pipe_out (39) = '1' or pipe_out (40) = '1' or pipe_out (41) = '1' or pipe_out (42) = '1' or pipe_out (43) = '1' or pipe_out (44) = '1' or pipe_out (45) = '1' or pipe_out (46) = '1' or pipe_out (47) = '1' or pipe_out (48) = '1' or pipe_out (49) = '1' or pipe_out (50) = '1' or pipe_out (51) = '1' or pipe_out (52) = '1' or pipe_out (53) = '1' or pipe_out (54) = '1' or pipe_out (55) = '1' or pipe_out (56) = '1' or pipe_out (57) = '1' or pipe_out (58) = '1' or pipe_out (59) = '1' or pipe_out (60) = '1' or pipe_out (61) = '1' or pipe_out (62) = '1' or pipe_out (63) = '1' or pipe_out (64) = '1' or pipe_out (65) = '1' or pipe_out (66) = '1' or pipe_out (67) = '1' or pipe_out (68) = '1' or pipe_out (69) = '1' or pipe_out (70) = '1' or pipe_out (71) = '1' or pipe_out (72) = '1' or pipe_out (73) = '1' or pipe_out (74) = '1' or pipe_out (75) = '1' or pipe_out (76) = '1' or pipe_out (77) = '1' or pipe_out (78) = '1' or pipe_out (79) = '1' or pipe_out (80) = '1' or pipe_out (81) = '1' or pipe_out (82) = '1' or pipe_out (83) = '1' or pipe_out (84) = '1' or pipe_out (85) = '1' or pipe_out (86) = '1' or pipe_out (87) = '1' or pipe_out (88) = '1' or pipe_out (89) = '1' or pipe_out (90) = '1' or pipe_out (91) = '1' or pipe_out (92) = '1' or pipe_out (93) = '1' or pipe_out (94) = '1' or pipe_out (95) = '1' or pipe_out (96) = '1' or pipe_out (97) = '1' or pipe_out (98) = '1' or (false) else '0';
pipe_in (99) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (100) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (101) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (102) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (103) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (104) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (105) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (106) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (107) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (108) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (109) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (3) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (110) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (111) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (112) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (113) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (114) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (115) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (116) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (117) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (118) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (119) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (120) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (121) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (122) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (123) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (124) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (125) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (126) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (127) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (128) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (129) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (130) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (131) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (132) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (133) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (134) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (135) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (136) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (137) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (138) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (139) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (140) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (141) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (142) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (143) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (144) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (145) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (146) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (147) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (148) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and (true) else '0';
pipe_in (149) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (150) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and (true) else '0';
pipe_in (151) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (152) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and (true) else '0';
pipe_in (153) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (154) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (155) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (156) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (157) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (158) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (159) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (160) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (161) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (162) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (163) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (164) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (0) = '1' and (true) else '0';
dataout (1) <= '1' when pipe_out (99) = '1' or pipe_out (100) = '1' or pipe_out (101) = '1' or pipe_out (102) = '1' or pipe_out (103) = '1' or pipe_out (104) = '1' or pipe_out (105) = '1' or pipe_out (106) = '1' or pipe_out (107) = '1' or pipe_out (108) = '1' or pipe_out (109) = '1' or pipe_out (110) = '1' or pipe_out (111) = '1' or pipe_out (112) = '1' or pipe_out (113) = '1' or pipe_out (114) = '1' or pipe_out (115) = '1' or pipe_out (116) = '1' or pipe_out (117) = '1' or pipe_out (118) = '1' or pipe_out (119) = '1' or pipe_out (120) = '1' or pipe_out (121) = '1' or pipe_out (122) = '1' or pipe_out (123) = '1' or pipe_out (124) = '1' or pipe_out (125) = '1' or pipe_out (126) = '1' or pipe_out (127) = '1' or pipe_out (128) = '1' or pipe_out (129) = '1' or pipe_out (130) = '1' or pipe_out (131) = '1' or pipe_out (132) = '1' or pipe_out (133) = '1' or pipe_out (134) = '1' or pipe_out (135) = '1' or pipe_out (136) = '1' or pipe_out (137) = '1' or pipe_out (138) = '1' or pipe_out (139) = '1' or pipe_out (140) = '1' or pipe_out (141) = '1' or pipe_out (142) = '1' or pipe_out (143) = '1' or pipe_out (144) = '1' or pipe_out (145) = '1' or pipe_out (146) = '1' or pipe_out (147) = '1' or pipe_out (148) = '1' or pipe_out (149) = '1' or pipe_out (150) = '1' or pipe_out (151) = '1' or pipe_out (152) = '1' or pipe_out (153) = '1' or pipe_out (154) = '1' or pipe_out (155) = '1' or pipe_out (156) = '1' or pipe_out (157) = '1' or pipe_out (158) = '1' or pipe_out (159) = '1' or pipe_out (160) = '1' or pipe_out (161) = '1' or pipe_out (162) = '1' or pipe_out (163) = '1' or pipe_out (164) = '1' or (false) else '0';
pipe_in (165) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (166) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (167) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (168) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (169) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (170) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (171) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (4) = '1' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (172) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (173) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (174) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (175) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (176) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (177) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (178) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (179) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (180) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (181) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (182) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (183) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (184) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '1' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (185) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (186) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (187) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (188) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (189) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (190) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (191) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (7) = '1' and datain (6) = '1' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (192) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (193) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (194) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (195) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (196) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (197) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (198) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (199) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (200) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (201) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (202) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '1' and datain (4) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (203) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (204) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (205) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (206) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (207) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (208) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (209) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and (true) else '0';
pipe_in (210) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '1' and (true) else '0';
pipe_in (211) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (212) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and (true) else '0';
dataout (2) <= '1' when pipe_out (165) = '1' or pipe_out (166) = '1' or pipe_out (167) = '1' or pipe_out (168) = '1' or pipe_out (169) = '1' or pipe_out (170) = '1' or pipe_out (171) = '1' or pipe_out (172) = '1' or pipe_out (173) = '1' or pipe_out (174) = '1' or pipe_out (175) = '1' or pipe_out (176) = '1' or pipe_out (177) = '1' or pipe_out (178) = '1' or pipe_out (179) = '1' or pipe_out (180) = '1' or pipe_out (181) = '1' or pipe_out (182) = '1' or pipe_out (183) = '1' or pipe_out (184) = '1' or pipe_out (185) = '1' or pipe_out (186) = '1' or pipe_out (187) = '1' or pipe_out (188) = '1' or pipe_out (189) = '1' or pipe_out (190) = '1' or pipe_out (191) = '1' or pipe_out (192) = '1' or pipe_out (193) = '1' or pipe_out (194) = '1' or pipe_out (195) = '1' or pipe_out (196) = '1' or pipe_out (197) = '1' or pipe_out (198) = '1' or pipe_out (199) = '1' or pipe_out (200) = '1' or pipe_out (201) = '1' or pipe_out (202) = '1' or pipe_out (203) = '1' or pipe_out (204) = '1' or pipe_out (205) = '1' or pipe_out (206) = '1' or pipe_out (207) = '1' or pipe_out (208) = '1' or pipe_out (209) = '1' or pipe_out (210) = '1' or pipe_out (211) = '1' or pipe_out (212) = '1' or (false) else '0';
pipe_in (213) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (214) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (215) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (216) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (217) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (1) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (218) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (219) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (220) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (221) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (222) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (3) = '1' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (223) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (224) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (225) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (226) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (227) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (228) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (229) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (230) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (231) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (232) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (233) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (5) = '1' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (234) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (235) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (236) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '1' and datain (4) = '1' and (true) else '0';
pipe_in (237) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (238) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '0' and (true) else '0';
pipe_in (239) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (2) = '1' and datain (1) = '0' and (true) else '0';
pipe_in (240) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (3) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (241) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (242) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (243) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (244) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (5) = '1' and datain (4) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (245) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and (true) else '0';
pipe_in (246) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '1' and datain (7) = '0' and datain (5) = '0' and (true) else '0';
pipe_in (247) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '1' and (true) else '0';
pipe_in (248) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '1' and (true) else '0';
pipe_in (249) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (250) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (251) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (252) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (253) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (254) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and (true) else '0';
dataout (3) <= '1' when pipe_out (213) = '1' or pipe_out (214) = '1' or pipe_out (215) = '1' or pipe_out (216) = '1' or pipe_out (217) = '1' or pipe_out (218) = '1' or pipe_out (219) = '1' or pipe_out (220) = '1' or pipe_out (221) = '1' or pipe_out (222) = '1' or pipe_out (223) = '1' or pipe_out (224) = '1' or pipe_out (225) = '1' or pipe_out (226) = '1' or pipe_out (227) = '1' or pipe_out (228) = '1' or pipe_out (229) = '1' or pipe_out (230) = '1' or pipe_out (231) = '1' or pipe_out (232) = '1' or pipe_out (233) = '1' or pipe_out (234) = '1' or pipe_out (235) = '1' or pipe_out (236) = '1' or pipe_out (237) = '1' or pipe_out (238) = '1' or pipe_out (239) = '1' or pipe_out (240) = '1' or pipe_out (241) = '1' or pipe_out (242) = '1' or pipe_out (243) = '1' or pipe_out (244) = '1' or pipe_out (245) = '1' or pipe_out (246) = '1' or pipe_out (247) = '1' or pipe_out (248) = '1' or pipe_out (249) = '1' or pipe_out (250) = '1' or pipe_out (251) = '1' or pipe_out (252) = '1' or pipe_out (253) = '1' or pipe_out (254) = '1' or (false) else '0';
pipe_in (255) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and datain (1) = '1' and datain (0) = '1' and (true) else '0';
pipe_in (256) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (6) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '1' and datain (0) = '0' and (true) else '0';
pipe_in (257) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '1' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (258) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (259) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (260) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (261) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '1' and datain (4) = '0' and datain (3) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (262) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (4) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (263) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (264) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (265) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '1' and datain (8) = '0' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (266) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (0) = '0' and (true) else '0';
pipe_in (267) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (268) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (269) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '1' and datain (6) = '1' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (270) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (271) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '1' and datain (5) = '1' and (true) else '0';
pipe_in (272) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '1' and datain (5) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (273) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and (true) else '0';
pipe_in (274) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (275) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (276) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (277) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '1' and (true) else '0';
pipe_in (278) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and (true) else '0';
dataout (4) <= '1' when pipe_out (255) = '1' or pipe_out (256) = '1' or pipe_out (257) = '1' or pipe_out (258) = '1' or pipe_out (259) = '1' or pipe_out (260) = '1' or pipe_out (261) = '1' or pipe_out (262) = '1' or pipe_out (263) = '1' or pipe_out (264) = '1' or pipe_out (265) = '1' or pipe_out (266) = '1' or pipe_out (267) = '1' or pipe_out (268) = '1' or pipe_out (269) = '1' or pipe_out (270) = '1' or pipe_out (271) = '1' or pipe_out (272) = '1' or pipe_out (273) = '1' or pipe_out (274) = '1' or pipe_out (275) = '1' or pipe_out (276) = '1' or pipe_out (277) = '1' or pipe_out (278) = '1' or (false) else '0';
pipe_in (279) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '1' and datain (2) = '0' and datain (1) = '0' and (true) else '0';
pipe_in (280) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (1) = '1' and (true) else '0';
pipe_in (281) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and datain (2) = '1' and (true) else '0';
pipe_in (282) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '1' and datain (3) = '1' and (true) else '0';
pipe_in (283) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (6) = '1' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and (true) else '0';
pipe_in (284) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (285) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '1' and (true) else '0';
pipe_in (286) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (3) = '0' and (true) else '0';
pipe_in (287) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '1' and datain (7) = '1' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and (true) else '0';
pipe_in (288) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (5) = '0' and datain (4) = '1' and datain (2) = '0' and (true) else '0';
pipe_in (289) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (6) = '0' and datain (5) = '0' and datain (2) = '1' and (true) else '0';
pipe_in (290) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (1) = '1' and (true) else '0';
pipe_in (291) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (0) = '1' and (true) else '0';
pipe_in (292) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (7) = '0' and datain (6) = '1' and (true) else '0';
pipe_in (293) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (6) = '0' and datain (5) = '1' and (true) else '0';
pipe_in (294) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '1' and (true) else '0';
dataout (5) <= '1' when pipe_out (279) = '1' or pipe_out (280) = '1' or pipe_out (281) = '1' or pipe_out (282) = '1' or pipe_out (283) = '1' or pipe_out (284) = '1' or pipe_out (285) = '1' or pipe_out (286) = '1' or pipe_out (287) = '1' or pipe_out (288) = '1' or pipe_out (289) = '1' or pipe_out (290) = '1' or pipe_out (291) = '1' or pipe_out (292) = '1' or pipe_out (293) = '1' or pipe_out (294) = '1' or (false) else '0';
pipe_in (295) <= '1' when datain (14) = '0' and datain (13) = '0' and datain (12) = '0' and datain (11) = '0' and datain (10) = '0' and datain (9) = '0' and datain (8) = '0' and datain (7) = '0' and datain (6) = '0' and datain (5) = '0' and datain (4) = '0' and datain (3) = '0' and datain (2) = '0' and datain (1) = '0' and datain (0) = '0' and (true) else '0';
dataout (6) <= '1' when pipe_out (295) = '1' or (false) else '0';
dataout (7) <= '0';

dataout (8) <= '0';

dataout (9) <= '0';

dataout (10) <= '0';

dataout (11) <= '0';

dataout (12) <= '0';

dataout (13) <= '0';

dataout (14) <= '0';


end Behavioural;
